LIBRARY IEEE ;
USE IEEE . STD_LOGIC_1164 . ALL ;
ENTITY AND_GATE IS
	PORT ( A , B : IN STD_LOGIC ;
		   F : OUT STD_LOGIC ) ;
END AND_GATE ;
ARCHITECTURE FUNC OF AND_GATE IS
BEGIN
	F <= A AND B ;
END FUNC ;
LIBRARY IEEE ;
USE IEEE . STD_LOGIC_1164 . ALL ;
ENTITY XOR_GATE IS
	PORT ( A , B : IN STD_LOGIC ;
		   F : OUT STD_LOGIC ) ;
END XOR_GATE ;
ARCHITECTURE FUNC OF XOR_GATE IS
BEGIN
	F <= A XOR B ;
END FUNC ;
LIBRARY IEEE ;
USE IEEE . STD_LOGIC_1164 . ALL ;
ENTITY HALF_ADDER IS
	PORT ( A , B : IN STD_LOGIC ;
	  SUM , COUT : OUT STD_LOGIC ) ;
END HALF_ADDER ;
ARCHITECTURE FUNC OF HALF_ADDER IS
	COMPONENT AND_GATE IS
		PORT ( A , B : IN STD_LOGIC ;
			   F : OUT STD_LOGIC ) ;
	END COMPONENT ;
	COMPONENT XOR_GATE IS
		PORT ( A , B : IN STD_LOGIC ;
			   F : OUT STD_LOGIC ) ;
	END COMPONENT ;
BEGIN
	G1 : XOR_GATE PORT MAP ( A , B , SUM ) ;
	G2 : AND_GATE PORT MAP ( A , B , COUT ) ;
END FUNC ;