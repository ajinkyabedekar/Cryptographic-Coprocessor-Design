LIBRARY IEEE ;
USE IEEE . STD_LOGIC_1164 . ALL ;
ENTITY NON_LINEAR_LOOKUP_TABLE IS
	PORT
	(
		LUTIN : IN STD_LOGIC_VECTOR ( 7 DOWNTO 0 ) ;
		LUTOUT : OUT STD_LOGIC_VECTOR ( 7 DOWNTO 0 )
	) ;
END NON_LINEAR_LOOKUP_TABLE ;
ARCHITECTURE FUNC OF NON_LINEAR_LOOKUP_TABLE IS
	SIGNAL MSN_IN , LSN_IN , MSN_OUT , LSN_OUT : STD_LOGIC_VECTOR ( 3 DOWNTO 0 ) ;
BEGIN
	MSN_IN <= LUTIN ( 7 DOWNTO 4 ) ;
	LSN_IN <= LUTIN ( 3 DOWNTO 0 ) ;
	SBOX_1 : PROCESS ( MSN_IN )
	BEGIN
		CASE ( MSN_IN ) IS
			WHEN "0000" => MSN_OUT <= "0001" ;
			WHEN "0001" => MSN_OUT <= "1011" ;
			WHEN "0010" => MSN_OUT <= "1001" ;
			WHEN "0011" => MSN_OUT <= "1100" ;
			WHEN "0100" => MSN_OUT <= "1101" ;
			WHEN "0101" => MSN_OUT <= "0110" ;
			WHEN "0110" => MSN_OUT <= "1111" ;
			WHEN "0111" => MSN_OUT <= "0011" ;
			WHEN "1000" => MSN_OUT <= "1110" ;
			WHEN "1001" => MSN_OUT <= "1000" ;
			WHEN "1010" => MSN_OUT <= "0111" ;
			WHEN "1011" => MSN_OUT <= "0100" ;
			WHEN "1100" => MSN_OUT <= "1010" ;
			WHEN "1101" => MSN_OUT <= "0010" ;
			WHEN "1110" => MSN_OUT <= "0101" ;
			WHEN "1111" => MSN_OUT <= "0000" ;
			WHEN OTHERS => MSN_OUT <= "0000" ;
		END CASE ;
	END PROCESS ;
	SBOX_2 : PROCESS ( LSN_IN )
	BEGIN
		CASE ( LSN_IN ) IS
			WHEN "0000" => LSN_OUT <= "1111" ;
			WHEN "0001" => LSN_OUT <= "0000" ;
			WHEN "0010" => LSN_OUT <= "1101" ;
			WHEN "0011" => LSN_OUT <= "0111" ;
			WHEN "0100" => LSN_OUT <= "1011" ;
			WHEN "0101" => LSN_OUT <= "1110" ;
			WHEN "0110" => LSN_OUT <= "0101" ;
			WHEN "0111" => LSN_OUT <= "1010" ;
			WHEN "1000" => LSN_OUT <= "1001" ;
			WHEN "1001" => LSN_OUT <= "0010" ;
			WHEN "1010" => LSN_OUT <= "1100" ;
			WHEN "1011" => LSN_OUT <= "0001" ;
			WHEN "1100" => LSN_OUT <= "0011" ;
			WHEN "1101" => LSN_OUT <= "0100" ;
			WHEN "1110" => LSN_OUT <= "1000" ;
			WHEN "1111" => LSN_OUT <= "0110" ;
			WHEN OTHERS => LSN_OUT <= "0000" ;
		END CASE ;
	END PROCESS ;
	LUTOUT <= MSN_OUT & LSN_OUT ;
END FUNC ;