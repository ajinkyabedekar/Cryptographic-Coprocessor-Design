LIBRARY IEEE ;
USE IEEE . STD_LOGIC_1164 . ALL ;
ENTITY AND_GATE IS
	PORT
	(
		A , B : IN STD_LOGIC ;
		    F : OUT STD_LOGIC
	) ;
END AND_GATE ;
ARCHITECTURE FUNC OF AND_GATE IS
BEGIN
	F <= A AND B ;
END FUNC ;

LIBRARY IEEE ;
USE IEEE . STD_LOGIC_1164 . ALL ;
ENTITY NOT_GATE IS
	PORT
	(
		A : IN STD_LOGIC ;
		F : OUT STD_LOGIC
	) ;
END NOT_GATE ;
ARCHITECTURE FUNC OF NOT_GATE IS
BEGIN
	F <= NOT A ;
END FUNC ;

LIBRARY IEEE ;
USE IEEE . STD_LOGIC_1164 . ALL ;
ENTITY ONE_TO_TWO_MUX_USING_AND_OR_NOT IS
	PORT
	(
		F , X : IN STD_LOGIC ;
		A , B : OUT STD_LOGIC
	) ;
END ONE_TO_TWO_MUX_USING_AND_OR_NOT ;
ARCHITECTURE FUNC OF ONE_TO_TWO_MUX_USING_AND_OR_NOT IS
	SIGNAL NOT_TO_AND : STD_LOGIC ;
BEGIN
	G1 : ENTITY WORK . NOT_GATE PORT MAP ( X , NOT_TO_AND ) ;
	G2 : ENTITY WORK . AND_GATE PORT MAP ( NOT_TO_AND , F , A ) ;
	G3 : ENTITY WORK . AND_GATE PORT MAP ( F , X , B ) ;
END FUNC ;