LIBRARY IEEE ;
USE IEEE . STD_LOGIC_1164 . ALL ;
ENTITY FULL_ADDER IS
	PORT
	(
		X , Y , C_IN : IN STD_LOGIC ;
		S , C_OUT : OUT STD_LOGIC
	) ;
END FULL_ADDER ;
ARCHITECTURE FUNC OF FULL_ADDER IS
BEGIN
	S <= X XOR Y XOR C_IN ;
	C_OUT <= ( X AND Y ) OR ( Y AND C_IN ) OR ( X AND C_IN ) ;
END FUNC ;