LIBRARY IEEE ;
USE IEEE . STD_LOGIC_1164 . ALL ;
ENTITY TWO_BIT_COMPARATOR IS
	PORT
	(
		A , B : IN STD_LOGIC_VECTOR ( 1 DOWNTO 0 ) ;
		A_LESS_THAN_B , A_EQUAL_TO_B , A_GREATER_THAN_B : OUT STD_LOGIC
	) ;
END TWO_BIT_COMPARATOR ;
ARCHITECTURE FUNC OF TWO_BIT_COMPARATOR IS
	SIGNAL TEMP1 , TEMP2 , TEMP3 , TEMP4 , TEMP5 , TEMP6 , TEMP7 , TEMP8 : STD_LOGIC ;
BEGIN
	TEMP1 <= A ( 1 ) XNOR B ( 1 ) ;
	TEMP2 <= A ( 0 ) XNOR B ( 0 ) ;
	A_EQUAL_TO_B <= TEMP1 AND TEMP2 ;
	TEMP3 <= ( NOT A ( 0 ) ) AND ( NOT A ( 1 ) ) AND B ( 0 ) ;
	TEMP4 <= ( NOT A ( 1 ) ) AND B ( 1 ) ;
	TEMP5 <= ( NOT A ( 0 ) ) AND B ( 1 ) AND B ( 0 ) ;
	A_LESS_THAN_B <= TEMP3 OR TEMP4 OR TEMP5 ;
	TEMP6 <= ( NOT B ( 0 ) ) AND ( NOT B ( 1 ) ) AND A ( 0 ) ;
	TEMP7 <= ( NOT B ( 1 ) ) AND A ( 1 ) ;
	TEMP8 <= ( NOT B ( 0 ) ) AND A ( 1 ) AND A ( 0 ) ;
	A_GREATER_THAN_B <= TEMP6 OR TEMP7 OR TEMP8 ;
END FUNC ;