LIBRARY IEEE ;
USE IEEE . STD_LOGIC_1164 . ALL ;
ENTITY NAND_GATE IS
	PORT ( A , B : IN STD_LOGIC ;
		   F : OUT STD_LOGIC ) ;
END NAND_GATE ;
ARCHITECTURE FUNC OF NAND_GATE IS
BEGIN
	F <= A NAND B ;
END FUNC ;