LIBRARY IEEE ;
USE IEEE . STD_LOGIC_1164 . ALL ;
ENTITY XNOR_GATE IS
	PORT ( A , B : IN STD_LOGIC ;
		   F : OUT STD_LOGIC ) ;
END XNOR_GATE ;
ARCHITECTURE FUNC OF XNOR_GATE IS
BEGIN
	F <= A XNOR B ;
END FUNC ;