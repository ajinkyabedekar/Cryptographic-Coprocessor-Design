LIBRARY IEEE ;
USE IEEE . STD_LOGIC_1164 . ALL ;
USE IEEE . STD_LOGIC_UNSIGNED . ALL ;
ENTITY TRAFFIC_LIGHT_CONTROLLER IS
	PORT
	(
		SENSOR , CLK , RESET : IN STD_LOGIC ;
		LIGHT_HIGHWAY , LIGHT_FARM : OUT STD_LOGIC_VECTOR ( 2 DOWNTO 0 )
	) ;
END TRAFFIC_LIGHT_CONTROLLER ;
ARCHITECTURE FUNC OF TRAFFIC_LIGHT_CONTROLLER IS
	SIGNAL COUNTER : STD_LOGIC_VECTOR ( 27 DOWNTO 0 ) := X"0000000" ;
	SIGNAL DELAY_COUNT : STD_LOGIC_VECTOR ( 3 DOWNTO 0 ) := X"0" ;
	SIGNAL DELAY_10_S , DELAY_3_S_FARM , DELAY_3_S_HIGHWAY , RED_LIGHT_ENABLE , YELLOW_LIGHT_1_ENABLE , YELLOW_LIGHT_2_ENABLE : STD_LOGIC := '0' ;
	SIGNAL CLK_ENABLE : STD_LOGIC ;
	TYPE FSM_STATES IS ( HIGHWAY_GREEN_FARM_RED , HIGHWAY_YELLOW_FARM_RED , HIGHWAY_RED_FARM_GREEN , HIGHWAY_RED_FARM_YELLOW ) ;
	SIGNAL CURRENT_STATE , NEXT_STATE : FSM_STATES ;
BEGIN
	PROCESS ( CLK , RESET )
	BEGIN
		IF ( RESET = '0' ) THEN
			CURRENT_STATE <= HIGHWAY_GREEN_FARM_RED ;
		ELSIF ( RISING_EDGE ( CLK ) ) THEN
			CURRENT_STATE <= NEXT_STATE ;
		END IF ;
	END PROCESS ;
	PROCESS ( CURRENT_STATE , SENSOR , DELAY_3_S_FARM , DELAY_3_S_HIGHWAY , DELAY_10_S )
	BEGIN
		CASE CURRENT_STATE IS
			WHEN HIGHWAY_GREEN_FARM_RED =>
				RED_LIGHT_ENABLE <= '0' ;
				YELLOW_LIGHT_1_ENABLE <= '0' ;
				YELLOW_LIGHT_2_ENABLE <= '0' ;
				LIGHT_HIGHWAY <= "001" ;
				LIGHT_FARM <= "100" ;
				IF ( SENSOR = '1' ) THEN
					NEXT_STATE <= HIGHWAY_YELLOW_FARM_RED ;
				ELSE
					NEXT_STATE <= HIGHWAY_GREEN_FARM_RED ;
				END IF ;
			WHEN HIGHWAY_YELLOW_FARM_RED =>
				LIGHT_HIGHWAY <= "010" ;
				LIGHT_FARM <= "100" ;
				RED_LIGHT_ENABLE <= '0' ;
				YELLOW_LIGHT_1_ENABLE <= '1' ;
				YELLOW_LIGHT_2_ENABLE <= '0' ;
				IF ( DELAY_3_S_HIGHWAY = '1' ) THEN
					NEXT_STATE <= HIGHWAY_RED_FARM_GREEN ;
				ELSE
					NEXT_STATE <= HIGHWAY_YELLOW_FARM_RED ;
				END IF ;
			WHEN HIGHWAY_RED_FARM_GREEN =>
				LIGHT_HIGHWAY <= "100" ;
				LIGHT_FARM <= "001" ;
				RED_LIGHT_ENABLE <= '1' ;
				YELLOW_LIGHT_1_ENABLE <= '0' ;
				YELLOW_LIGHT_2_ENABLE <= '0' ;
				IF ( DELAY_10_S = '1' ) THEN
					NEXT_STATE <= HIGHWAY_RED_FARM_YELLOW ;
				ELSE
					NEXT_STATE <= HIGHWAY_RED_FARM_GREEN ;
				END IF ;
			WHEN HIGHWAY_RED_FARM_YELLOW =>
				LIGHT_HIGHWAY <= "100" ;
				LIGHT_FARM <= "010" ;
				RED_LIGHT_ENABLE <= '0' ;
				YELLOW_LIGHT_1_ENABLE <= '0' ;
				YELLOW_LIGHT_2_ENABLE <= '1' ;
				IF ( DELAY_3_S_FARM = '1' ) THEN
					NEXT_STATE <= HIGHWAY_GREEN_FARM_RED ;
				ELSE
					NEXT_STATE <= HIGHWAY_RED_FARM_YELLOW ;
				END IF ;
			WHEN OTHERS => NEXT_STATE <= HIGHWAY_GREEN_FARM_RED ;
		END CASE ;
	END PROCESS ;
	PROCESS ( CLK )
	BEGIN
		IF ( RISING_EDGE ( CLK ) ) THEN
			IF ( CLK_ENABLE = '1' ) THEN
				IF ( RED_LIGHT_ENABLE = '1' OR YELLOW_LIGHT_1_ENABLE = '1' OR YELLOW_LIGHT_2_ENABLE = '1' ) THEN
					DELAY_COUNT <= DELAY_COUNT + X"1" ;
					IF ( ( DELAY_COUNT = X"9" ) AND RED_LIGHT_ENABLE = '1' ) THEN
						DELAY_10_S <= '1' ;
						DELAY_3_S_HIGHWAY <= '0' ;
						DELAY_3_S_FARM <= '0' ;
						DELAY_COUNT <= X"0" ;
					ELSIF ( ( DELAY_COUNT = X"2" ) AND YELLOW_LIGHT_1_ENABLE = '1' ) THEN
						DELAY_10_S <= '0' ;
						DELAY_3_S_HIGHWAY <= '1' ;
						DELAY_3_S_FARM <= '0' ;
						DELAY_COUNT <= X"0" ;
					ELSIF ( ( DELAY_COUNT = X"2" ) AND YELLOW_LIGHT_2_ENABLE = '1' ) THEN
						DELAY_10_S <= '0' ;
						DELAY_3_S_HIGHWAY <= '0' ;
						DELAY_3_S_FARM <= '1' ;
						DELAY_COUNT <= X"0" ;
					ELSE
						DELAY_10_S <= '0' ;
						DELAY_3_S_HIGHWAY <= '0' ;
						DELAY_3_S_FARM <= '0' ;
					END IF ;
				END IF ;
			END IF ;
		END IF ;
	END PROCESS ;
	PROCESS ( CLK )
	BEGIN
		IF ( RISING_EDGE ( CLK ) ) THEN
			COUNTER <= COUNTER + X"0000001" ;
			IF ( COUNTER >= X"0000003" ) THEN
				COUNTER <= X"0000000" ;
			END IF ;
		END IF ;
	END PROCESS ;
	CLK_ENABLE <= '1' WHEN COUNTER = X"0003" ELSE '0' ;
END FUNC ;