LIBRARY IEEE ;
USE IEEE . STD_LOGIC_1164 . ALL ;
ENTITY COMBINATIONAL_LOGIC_UNIT_OF_COPROCESSOR IS
	PORT
	(
		A_BUS : IN STD_LOGIC_VECTOR ( 15 DOWNTO 0 ) ;
		B_BUS : IN STD_LOGIC_VECTOR ( 15 DOWNTO 0 ) ;
		CTRL : IN STD_LOGIC_VECTOR ( 3 DOWNTO 0 ) ;
		RESULT : OUT STD_LOGIC_VECTOR ( 15 DOWNTO 0 )
	) ;
END COMBINATIONAL_LOGIC_UNIT_OF_COPROCESSOR ;
ARCHITECTURE FUNC OF COMBINATIONAL_LOGIC_UNIT_OF_COPROCESSOR IS
	COMPONENT NON_LINEAR_LOOKUP_TABLE IS
	PORT
	(
		LUTIN : IN STD_LOGIC_VECTOR ( 7 DOWNTO 0 ) ;
		LUTOUT : OUT STD_LOGIC_VECTOR ( 7 DOWNTO 0 )
	) ;
	END COMPONENT NON_LINEAR_LOOKUP_TABLE ;
	COMPONENT SHIFTER IS
	GENERIC
	(
		N : INTEGER := 16
	) ;
	PORT
	(
		SHIFT_INPUT : IN STD_LOGIC_VECTOR ( N - 1 DOWNTO 0 ) ;
		SHIFT_CTRL : IN STD_LOGIC_VECTOR ( 3 DOWNTO 0 ) ;
		SHIFT_OUT : OUT STD_LOGIC_VECTOR ( N - 1 DOWNTO 0 )
	) ;
	END COMPONENT SHIFTER ;
	COMPONENT SIXTEEN_BIT_ALU IS
	PORT
	(
		ABUS : IN STD_LOGIC_VECTOR ( 15 DOWNTO 0 ) ;
		BBUS : IN STD_LOGIC_VECTOR ( 15 DOWNTO 0 ) ;
		ALUCTRL : IN STD_LOGIC_VECTOR ( 3 DOWNTO 0 ) ;
		ALUOUT : OUT STD_LOGIC_VECTOR ( 15 DOWNTO 0 )
	) ;
	END COMPONENT SIXTEEN_BIT_ALU ;
	SIGNAL TEMP_OUT_1 , TEMP_OUT_2 , TEMP_OUT_3 : STD_LOGIC_VECTOR ( 15 DOWNTO 0 ) ;
	SIGNAL LUT_OUT : STD_LOGIC_VECTOR ( 7 DOWNTO 0 ) ;
BEGIN
	ALU_UNIT : SIXTEEN_BIT_ALU PORT MAP ( ABUS => A_BUS , BBUS => B_BUS , ALUCTRL => CTRL , ALUOUT => TEMP_OUT_1 ) ;
	SHIFTER_UNIT : SHIFTER GENERIC MAP ( N => 16 )
	PORT MAP ( SHIFT_INPUT => B_BUS , SHIFT_CTRL => CTRL , SHIFT_OUT => TEMP_OUT_2 ) ;
	NON_LINEAR_LOOKUP_UNIT : NON_LINEAR_LOOKUP_TABLE
	PORT MAP ( LUTIN => A_BUS ( 7 DOWNTO 0 ) , LUTOUT => LUT_OUT ) ;
	TEMP_OUT_3 <= A_BUS ( 15 DOWNTO 8 ) & LUT_OUT ;
	CONTROL_LOGIC : PROCESS ( CTRL , TEMP_OUT_1 , TEMP_OUT_3 , TEMP_OUT_2 )
	BEGIN
		CASE ( CTRL ( 3 DOWNTO 3 ) ) IS
			WHEN "0" => RESULT <= TEMP_OUT_1 ;
			WHEN OTHERS =>
				CASE ( CTRL ( 1 DOWNTO 0 ) ) IS
					WHEN "11" => RESULT <= TEMP_OUT_3 ;
					WHEN OTHERS => RESULT <= TEMP_OUT_2 ;
				END CASE ;
		END CASE ;
	END PROCESS CONTROL_LOGIC ;
END FUNC;