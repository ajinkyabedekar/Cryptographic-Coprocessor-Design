LIBRARY IEEE ;
USE IEEE . STD_LOGIC_1164 . ALL ;
ENTITY N_BIT_ADDER IS
	PORT
	(
		INPUT_1 , INPUT_2 : IN STD_LOGIC_VECTOR ( 31 DOWNTO 0 ) ;
		ANSWER : OUT STD_LOGIC_VECTOR ( 31 DOWNTO 0 ) ;
		I_CLOCK : STD_LOGIC
	) ;
END N_BIT_ADDER ;
ARCHITECTURE FUNC OF N_BIT_ADDER IS
	COMPONENT HALF_ADDER IS
		PORT
		(
			X , Y : IN STD_LOGIC ;
			S , C : OUT STD_LOGIC
		) ;
	END COMPONENT ;
	COMPONENT FULL_ADDER IS
		PORT
		(
			X , Y , C_IN : IN STD_LOGIC ;
			S , C_OUT : OUT STD_LOGIC
		) ;
	END COMPONENT ;
	SIGNAL CARRY_OUT : STD_LOGIC ;
	SIGNAL CARRY : STD_LOGIC_VECTOR ( 31 DOWNTO 0 ) ;
BEGIN
	P1 : PROCESS ( I_CLOCK )
	BEGIN
		FOR II IN 0 TO 31 LOOP
			IF ( II = 0 ) THEN
				HALF_ADDER PORT MAP ( INPUT_1 ( 0 ) , INPUT_2 ( 0 ) , ANSWER ( 0 ) , CARRY ( 0 ) ) ;
			ELSE
				FULL_ADDER PORT MAP ( INPUT_1 ( II ) , INPUT_2 ( II ) , CARRY ( II - 1 ) , ANSWER ( II ) , CARRY ( II ) ) ;
			END IF ;
		END LOOP ;
		CARRY_OUT := CARRY ( 31 ) ;
	END PROCESS ;
END FUNC ;