LIBRARY IEEE ;
USE IEEE . STD_LOGIC_1164 . ALL ;
ENTITY ENCODER1 IS
	PORT (
	A : IN STD_LOGIC_VECTOR ( 3 DOWNTO 0 ) ;
	B : OUT STD_LOGIC_VECTOR ( 1 DOWNTO 0 )
	) ;
END ENCODER1 ;
ARCHITECTURE BHV OF ENCODER1 IS
BEGIN
PROCESS ( A )
BEGIN
	IF ( A = "1000" ) THEN
		B <= "00" ;
	ELSIF ( A = "0100" ) THEN
		B <= "01" ;
	ELSIF ( A = "0010" ) THEN
		B <= "10" ;
	ELSIF ( A = "0001" ) THEN
		B <= "11" ;
	ELSE
		B <= "ZZ" ;
	END IF ;
END PROCESS ;
END BHV ;




LIBRARY IEEE ;
USE IEEE . STD_LOGIC_1164 . ALL ;
ENTITY DECODER1 IS
	PORT (
	A : IN STD_LOGIC_VECTOR ( 1 DOWNTO 0 ) ;
	B : OUT STD_LOGIC_VECTOR ( 3 DOWNTO 0 )
	) ;
END DECODER1 ;
ARCHITECTURE BHV OF DECODER1 IS
BEGIN
PROCESS ( A )
BEGIN
	IF ( A = "00" ) THEN
		B <= "0001" ;
	ELSIF ( A = "01" ) THEN
		B <= "0010" ;
	ELSIF ( A = "10" ) THEN
		B <= "0100" ;
	ELSE
		B <= "1000" ;
	END IF ;
END PROCESS ;
END BHV ;