LIBRARY IEEE ;
USE IEEE . STD_LOGIC_1164 . ALL ;
ENTITY AND_GATE IS
	PORT ( A , B : IN STD_LOGIC ;
		   F : OUT STD_LOGIC ) ;
END AND_GATE ;
ARCHITECTURE FUNC OF AND_GATE IS
BEGIN
	F <= A AND B ;
END FUNC ;
LIBRARY IEEE ;
USE IEEE . STD_LOGIC_1164 . ALL ;
ENTITY OR_GATE IS
	PORT ( A , B : IN STD_LOGIC ;
		   F : OUT STD_LOGIC ) ;
END OR_GATE ;
ARCHITECTURE FUNC OF OR_GATE IS
BEGIN
	F <= A OR B ;
END FUNC ;
LIBRARY IEEE ;
USE IEEE . STD_LOGIC_1164 . ALL ;
ENTITY NOT_GATE IS
	PORT ( IN_PORT : IN STD_LOGIC ;
	      OUT_PORT : OUT STD_LOGIC ) ;
END NOT_GATE ;
ARCHITECTURE FUNC OF NOT_GATE IS
BEGIN
	OUT_PORT <= NOT IN_PORT ;
END FUNC ;
LIBRARY IEEE ;
USE IEEE . STD_LOGIC_1164 . ALL ;
ENTITY TWO_TO_ONE_MULTIPLEXER IS
	PORT ( D0 , D1 , S : IN STD_LOGIC ;
			 F : OUT STD_LOGIC ) ;
END TWO_TO_ONE_MULTIPLEXER ;
ARCHITECTURE FUNC OF TWO_TO_ONE_MULTIPLEXER IS
	COMPONENT AND_GATE IS
		PORT ( A , B : IN STD_LOGIC ;
			   F : OUT STD_LOGIC ) ;
	END COMPONENT ;
	COMPONENT OR_GATE IS
		PORT ( A , B : IN STD_LOGIC ;
			   F : OUT STD_LOGIC ) ;
	END COMPONENT ;
	COMPONENT NOT_GATE IS
		PORT ( IN_PORT : IN STD_LOGIC ;
		      OUT_PORT : OUT STD_LOGIC ) ;
	END COMPONENT ;
	SIGNAL AND_OUT_1 , AND_OUT_2 , INV_OUT : STD_LOGIC ;
BEGIN
	G1 : NOT_GATE PORT MAP ( S , INV_OUT ) ;
	G2 : AND_GATE PORT MAP ( INV_OUT , D0 , AND_OUT_1 ) ;
	G3 : AND_GATE PORT MAP ( S , D1 , AND_OUT_2 ) ;
	G4 : OR_GATE PORT MAP ( AND_OUT_1 , AND_OUT_2 , F ) ;
END FUNC ;




LIBRARY IEEE ;
USE IEEE . STD_LOGIC_1164 . ALL ;
ENTITY MUXUSINGWHEN IS
	PORT ( SEL : IN STD_LOGIC ;
		A : IN STD_LOGIC_VECTOR ( 3 DOWNTO 0 ) ;
		B : IN STD_LOGIC_VECTOR ( 3 DOWNTO 0 ) ;
		X : OUT STD_LOGIC_VECTOR ( 3 DOWNTO 0 ) ) ;
END MUXUSINGWHEN ;
ARCHITECTURE BEHAVIORAL OF MUXUSINGWHEN IS
BEGIN
	X <= A WHEN ( SEL = '1' ) ELSE B ;
END BEHAVIORAL ;




LIBRARY IEEE ;
USE IEEE . STD_LOGIC_1164 . ALL ;
ENTITY MUX_4TO1_TOP IS
	PORT ( SEL : IN STD_LOGIC_VECTOR ( 1 DOWNTO 0 ) ;
		A : STD_LOGIC_VECTOR ( 3 DOWNTO 0 ) ;
		X : OUT STD_LOGIC ) ;
END MUX_4TO1_TOP ;
ARCHITECTURE BEHAVIORAL OF MUX_4TO1_TOP IS
BEGIN
WITH SEL SELECT
	X <= A ( 0 ) WHEN "00" ,
		A (1) WHEN "01",
		A (2) WHEN "10",
		A (3) WHEN "11",
		'0' WHEN OTHERS;
END BEHAVIORAL ;