LIBRARY IEEE ;
USE IEEE . STD_LOGIC_1164 . ALL ;
ENTITY OR_GATE IS
	PORT
	(
		A , B : IN STD_LOGIC ;
		    F : OUT STD_LOGIC
	) ;
END OR_GATE ;
ARCHITECTURE FUNC OF OR_GATE IS
BEGIN
	F <= A OR B ;
END FUNC ;

LIBRARY IEEE ;
USE IEEE . STD_LOGIC_1164 . ALL ;
ENTITY NOT_GATE IS
	PORT
	(
		A : IN STD_LOGIC ;
		F : OUT STD_LOGIC
	) ;
END NOT_GATE ;
ARCHITECTURE FUNC OF NOT_GATE IS
BEGIN
	F <= NOT A ;
END FUNC ;

LIBRARY IEEE ;
USE IEEE . STD_LOGIC_1164 . ALL ;
ENTITY AND_GATE_USING_NOR_GATE IS
	PORT
	(
		A , B : IN STD_LOGIC ;
		    F : OUT STD_LOGIC
	) ;
END AND_GATE_USING_NOR_GATE ;
ARCHITECTURE FUNC OF AND_GATE_USING_NOR_GATE IS
	COMPONENT OR_GATE IS
		PORT
		(
			A , B : IN STD_LOGIC ;
			    F : OUT STD_LOGIC
		) ;
	END COMPONENT ;
	COMPONENT NOT_GATE IS
		PORT
		(
			A : IN STD_LOGIC ;
			F : OUT STD_LOGIC
		) ;
	END COMPONENT ;
	SIGNAL OR_TO_NOT_1 , OR_TO_NOT_2 , OR_TO_NOT_3 , NOT_TO_OR_1 , NOT_TO_OR_2 : STD_LOGIC ;
BEGIN
	G1 : OR_GATE PORT MAP ( A , A , OR_TO_NOT_1 ) ;
	G2 : NOT_GATE PORT MAP ( OR_TO_NOT_1 , NOT_TO_OR_1 ) ;
	G3 : OR_GATE PORT MAP ( B , B , OR_TO_NOT_2 ) ;
	G4 : NOT_GATE PORT MAP ( OR_TO_NOT_2 , NOT_TO_OR_2 ) ;
	G5 : OR_GATE PORT MAP ( NOT_TO_OR_1 , NOT_TO_OR_2 , OR_TO_NOT_3 ) ;
	G6 : NOT_GATE PORT MAP ( OR_TO_NOT_3 , F ) ;
END FUNC ;