LIBRARY IEEE ;
USE IEEE . STD_LOGIC_1164 . ALL ;
ENTITY HALF_ADDER IS
	PORT
	(
		X , Y : IN STD_LOGIC ;
		S , C : OUT STD_LOGIC
	) ;
END HALF_ADDER ;
ARCHITECTURE FUNC OF HALF_ADDER IS
BEGIN
	S <= X XOR Y ;
	C <= X AND Y ;
END FUNC ;