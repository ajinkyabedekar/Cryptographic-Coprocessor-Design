LIBRARY IEEE ;
USE IEEE . STD_LOGIC_1164 . ALL ;
ENTITY XOR_GATE IS
	PORT ( A , B : IN STD_LOGIC ;
		   F : OUT STD_LOGIC ) ;
END XOR_GATE ;
ARCHITECTURE FUNC OF XOR_GATE IS
BEGIN
	F <= A XOR B ;
END FUNC ;
LIBRARY IEEE ;
USE IEEE . STD_LOGIC_1164 . ALL ;
ENTITY FULL_ADDER IS
	PORT ( X , Y , CIN : IN STD_LOGIC ;
		SUM , COUT : OUT STD_LOGIC ) ;
END FULL_ADDER ;
ARCHITECTURE FUNC OF FULL_ADDER IS
BEGIN
	SUM <= ( X XOR Y ) XOR CIN ;
	COUT <= ( X AND ( Y OR CIN ) ) OR ( CIN AND Y ) ;
END FUNC ;
LIBRARY IEEE ;
USE IEEE . STD_LOGIC_1164 . ALL ;
ENTITY FOUR_BIT_ADDER_SUBTRACTOR IS
	PORT ( MODE : IN STD_LOGIC ;
  A3 , A2 , A1 , A0 : IN STD_LOGIC ;
  B3 , B2 , B1 , B0 : IN STD_LOGIC ;
  S3 , S2 , S1 , S0 : OUT STD_LOGIC ;
	   COUT , V : OUT STD_LOGIC ) ;
END FOUR_BIT_ADDER_SUBTRACTOR ;
ARCHITECTURE FUNC OF FOUR_BIT_ADDER_SUBTRACTOR IS
	COMPONENT XOR_GATE IS
		PORT ( A , B : IN STD_LOGIC ;
			   F : OUT STD_LOGIC ) ;
	END COMPONENT ;
	COMPONENT FULL_ADDER IS
		PORT ( X , Y , CIN : IN STD_LOGIC ;
			SUM , COUT : OUT STD_LOGIC ) ;
	END COMPONENT ;
	SIGNAL C1 , C2 , C3 , C4 : STD_LOGIC ;
	SIGNAL XOR_0 , XOR_1 , XOR_2 , XOR_3 : STD_LOGIC ;
BEGIN
	GX0 : XOR_GATE PORT MAP ( MODE , B0 , XOR_0 ) ;
	GX1 : XOR_GATE PORT MAP ( MODE , B1 , XOR_1 ) ;
	GX2 : XOR_GATE PORT MAP ( MODE , B2 , XOR_2 ) ;
	GX3 : XOR_GATE PORT MAP ( MODE , B3 , XOR_3 ) ;
	FA0 : FULL_ADDER PORT MAP ( A0 , XOR_0 , MODE , S0 , C1 ) ;
	FA1 : FULL_ADDER PORT MAP ( A1 , XOR_1 , C1 , S1 , C2 ) ;
	FA2 : FULL_ADDER PORT MAP ( A2 , XOR_2 , C2 , S2 , C3 ) ;
	FA3 : FULL_ADDER PORT MAP ( A3 , XOR_3 , C3 , S3 , C4 ) ;
	VOUT : XOR_GATE PORT MAP ( C3 , C4 , V ) ;
	COUT <= C4 ;
END FUNC ;