LIBRARY IEEE ;
USE IEEE . STD_LOGIC_1164 . ALL ;
ENTITY AND_GATE IS
	PORT
	(
		A , B : IN STD_LOGIC ;
		    F : OUT STD_LOGIC
	) ;
END AND_GATE ;
ARCHITECTURE FUNC OF AND_GATE IS
BEGIN
	F <= A AND B ;
END FUNC ;

LIBRARY IEEE ;
USE IEEE . STD_LOGIC_1164 . ALL ;
ENTITY OR_GATE IS
	PORT
	(
		A , B : IN STD_LOGIC ;
		    F : OUT STD_LOGIC
	) ;
END OR_GATE ;
ARCHITECTURE FUNC OF OR_GATE IS
BEGIN
	F <= A OR B ;
END FUNC ;

LIBRARY IEEE ;
USE IEEE . STD_LOGIC_1164 . ALL ;
ENTITY NOT_GATE IS
	PORT
	(
		A : IN STD_LOGIC ;
		F : OUT STD_LOGIC
	) ;
END NOT_GATE ;
ARCHITECTURE FUNC OF NOT_GATE IS
BEGIN
	F <= NOT A ;
END FUNC ;

LIBRARY IEEE ;
USE IEEE . STD_LOGIC_1164 . ALL ;
ENTITY TWO_TO_ONE_MUX_USING_AND_OR_NOT IS
	PORT
	(
		A , B , X : IN STD_LOGIC ;
			F : OUT STD_LOGIC
	) ;
END TWO_TO_ONE_MUX_USING_AND_OR_NOT ;
ARCHITECTURE FUNC OF TWO_TO_ONE_MUX_USING_AND_OR_NOT IS
	SIGNAL NOT_TO_AND , AND_TO_OR_1 , AND_TO_OR_2 : STD_LOGIC ;
BEGIN
	G1 : ENTITY WORK . NOT_GATE PORT MAP ( X , NOT_TO_AND ) ;
	G2 : ENTITY WORK . AND_GATE PORT MAP ( A , NOT_TO_AND , AND_TO_OR_1 ) ;
	G3 : ENTITY WORK . AND_GATE PORT MAP ( X , B , AND_TO_OR_2 ) ;
	G4 : ENTITY WORK . OR_GATE PORT MAP ( AND_TO_OR_1 , AND_TO_OR_2 , F ) ;
END FUNC ;

LIBRARY IEEE ;
USE IEEE . STD_LOGIC_1164 . ALL ;
ENTITY FOUR_TO_ONE_MUX_USING_TWO_TO_ONE_MUX IS
	PORT
	(
		A : IN STD_LOGIC_VECTOR ( 3 DOWNTO 0 ) ;
		S : IN STD_LOGIC_VECTOR ( 1 DOWNTO 0 ) ;
		F : OUT STD_LOGIC
	) ;
END FOUR_TO_ONE_MUX_USING_TWO_TO_ONE_MUX ;
ARCHITECTURE FUNC OF FOUR_TO_ONE_MUX_USING_TWO_TO_ONE_MUX IS
	SIGNAL MUX_TO_MUX_1 , MUX_TO_MUX_2 : STD_LOGIC ;
BEGIN
	G1 : ENTITY WORK . TWO_TO_ONE_MUX_USING_AND_OR_NOT PORT MAP ( A ( 0 ) , A ( 1 ) , S ( 0 ) , MUX_TO_MUX_1 ) ;
	G2 : ENTITY WORK . TWO_TO_ONE_MUX_USING_AND_OR_NOT PORT MAP ( A ( 2 ) , A ( 3 ) , S ( 0 ) , MUX_TO_MUX_2 ) ;
	G3 : ENTITY WORK . TWO_TO_ONE_MUX_USING_AND_OR_NOT PORT MAP ( MUX_TO_MUX_1 , MUX_TO_MUX_2 , S ( 1 ) , F ) ;
END FUNC ;