LIBRARY IEEE ;
USE IEEE . STD_LOGIC_1164 . ALL ;
ENTITY AND_GATE IS
	PORT
	(
		A , B : IN STD_LOGIC ;
		    F : OUT STD_LOGIC
	) ;
END AND_GATE ;
ARCHITECTURE FUNC OF AND_GATE IS
BEGIN
	F <= A AND B ;
END FUNC ;

LIBRARY IEEE ;
USE IEEE . STD_LOGIC_1164 . ALL ;
ENTITY NOT_GATE IS
	PORT
	(
		A : IN STD_LOGIC ;
		F : OUT STD_LOGIC
	) ;
END NOT_GATE ;
ARCHITECTURE FUNC OF NOT_GATE IS
BEGIN
	F <= NOT A ;
END FUNC ;

LIBRARY IEEE ;
USE IEEE . STD_LOGIC_1164 . ALL ;
ENTITY NAND_USING_AND_OR_NOT IS
	PORT
	(
		A , B : IN STD_LOGIC ;
		    F : OUT STD_LOGIC
	) ;
END NAND_USING_AND_OR_NOT ;
ARCHITECTURE FUNC OF NAND_USING_AND_OR_NOT IS
	COMPONENT AND_GATE IS
		PORT
		(
			A , B : IN STD_LOGIC ;
			    F : OUT STD_LOGIC
		) ;
	END COMPONENT ;
	COMPONENT NOT_GATE IS
		PORT
		(
			A : IN STD_LOGIC ;
			F : OUT STD_LOGIC
		) ;
	END COMPONENT ;
	SIGNAL AND_TO_NOT : STD_LOGIC ;
BEGIN
	G1 : AND_GATE PORT MAP ( A , B , AND_TO_NOT ) ;
	G2 : NOT_GATE PORT MAP ( AND_TO_NOT , F ) ;
END FUNC ;