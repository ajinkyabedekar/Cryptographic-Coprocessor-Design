LIBRARY IEEE ;
USE IEEE . STD_LOGIC_1164 . ALL ;
ENTITY SIXTEEN_BIT_ALU IS
	PORT
	(
		ABUS : IN STD_LOGIC_VECTOR ( 15 DOWNTO 0 ) ;
		BBUS : IN STD_LOGIC_VECTOR ( 15 DOWNTO 0 ) ;
		ALUCTRL : IN STD_LOGIC_VECTOR ( 3 DOWNTO 0 ) ;
		ALUOUT : OUT STD_LOGIC_VECTOR ( 15 DOWNTO 0 )
	) ;
END SIXTEEN_BIT_ALU ;
ARCHITECTURE FUNC OF SIXTEEN_BIT_ALU IS
	COMPONENT N_BIT_ADDER IS
		GENERIC
		(
			N : INTEGER := 32
		) ;
		PORT
		(
			INPUT_1 : IN STD_LOGIC_VECTOR ( N - 1 DOWNTO 0 ) ;
			INPUT_2 : IN STD_LOGIC_VECTOR ( N - 1 DOWNTO 0 ) ;
			ANSWER : OUT STD_LOGIC_VECTOR ( N - 1 DOWNTO 0 )
		) ;
	END COMPONENT N_BIT_ADDER ;
	SIGNAL BBUS_NOT : STD_LOGIC_VECTOR ( 16 - 1 DOWNTO 0 ) ;
	SIGNAL TEMP_OUT_1 : STD_LOGIC_VECTOR ( 16 - 1 DOWNTO 0 ) ;
	SIGNAL TEMP_OUT_2 : STD_LOGIC_VECTOR ( 16 - 1 DOWNTO 0 ) ;
	SIGNAL TEMP : STD_LOGIC_VECTOR ( 16 - 1 DOWNTO 0 ) ;
BEGIN
	U1_N_BIT_ADDER : N_BIT_ADDER GENERIC MAP ( N => 16 )
	PORT MAP ( INPUT_1 => ABUS , INPUT_2 => BBUS , ANSWER => TEMP_OUT_1 ) ;
	U2_N_BIT_ADDER : N_BIT_ADDER GENERIC MAP ( N => 16 )
	PORT MAP ( INPUT_1 => ABUS , INPUT_2 => BBUS_NOT , ANSWER => TEMP_OUT_2 ) ;
	U3_N_BIT_ADDER : N_BIT_ADDER GENERIC MAP ( N => 16 )
	PORT MAP ( INPUT_1 => TEMP_OUT_2 , INPUT_2 => x"0001" , ANSWER => TEMP ) ;
	BBUS_NOT <= NOT BBUS ;
	PROCESS ( ALUCTRL , ABUS , BBUS , TEMP_OUT_1 , TEMP )
	BEGIN
		CASE ( ALUCTRL ) IS
			WHEN "0000" =>  ALUOUT <= TEMP_OUT_1 ;
			WHEN "0001" =>  ALUOUT <= TEMP ;
			WHEN "0010" =>  ALUOUT <= ABUS AND BBUS ;
			WHEN "0011" =>  ALUOUT <= ABUS OR BBUS ;
			WHEN "0100" =>  ALUOUT <= ABUS XOR BBUS ;
			WHEN "0101" =>  ALUOUT <= NOT ABUS ;
			WHEN "0110" =>  ALUOUT <= ABUS ;
			WHEN OTHERS => ALUOUT <= TEMP_OUT_1 ;
		END CASE ;
	END PROCESS ;
END FUNC ;