LIBRARY IEEE ;
USE IEEE . STD_LOGIC_1164 . ALL ;
ENTITY AND_GATE IS
	PORT
	(
		A , B : IN STD_LOGIC ;
		    F : OUT STD_LOGIC
	) ;
END AND_GATE ;
ARCHITECTURE FUNC OF AND_GATE IS
BEGIN
	F <= A AND B ;
END FUNC ;

LIBRARY IEEE ;
USE IEEE . STD_LOGIC_1164 . ALL ;
ENTITY NOT_GATE IS
	PORT
	(
		A : IN STD_LOGIC ;
		F : OUT STD_LOGIC
	) ;
END NOT_GATE ;
ARCHITECTURE FUNC OF NOT_GATE IS
BEGIN
	F <= NOT A ;
END FUNC ;

LIBRARY IEEE ;
USE IEEE . STD_LOGIC_1164 . ALL ;
ENTITY XOR_GATE_USING_NAND_GATE IS
	PORT
	(
		A , B : IN STD_LOGIC ;
		    F : OUT STD_LOGIC
	) ;
END XOR_GATE_USING_NAND_GATE ;
ARCHITECTURE FUNC OF XOR_GATE_USING_NAND_GATE IS
	COMPONENT AND_GATE IS
		PORT
		(
			A , B : IN STD_LOGIC ;
			    F : OUT STD_LOGIC
		) ;
	END COMPONENT ;
	COMPONENT NOT_GATE IS
		PORT
		(
			A : IN STD_LOGIC ;
			F : OUT STD_LOGIC
		) ;
	END COMPONENT ;
	SIGNAL AND_TO_NOT_1 , AND_TO_NOT_2 , AND_TO_NOT_3 , AND_TO_NOT_4 , NOT_TO_AND_1 , NOT_TO_AND_2 , NOT_TO_AND_3 : STD_LOGIC ;
BEGIN
	G1 : AND_GATE PORT MAP ( A , B , AND_TO_NOT_1 ) ;
	G2 : NOT_GATE PORT MAP ( AND_TO_NOT_1 , NOT_TO_AND_1 ) ;
	G3 : AND_GATE PORT MAP ( A , NOT_TO_AND_1 , AND_TO_NOT_2 ) ;
	G4 : NOT_GATE PORT MAP ( AND_TO_NOT_2 , NOT_TO_AND_2 ) ;
	G5 : AND_GATE PORT MAP ( B , NOT_TO_AND_1 , AND_TO_NOT_3 ) ;
	G6 : NOT_GATE PORT MAP ( AND_TO_NOT_3 , NOT_TO_AND_3 ) ;
	G7 : AND_GATE PORT MAP ( NOT_TO_AND_2 , NOT_TO_AND_3 , AND_TO_NOT_4 ) ;
	G8 : NOT_GATE PORT MAP ( AND_TO_NOT_4 , F ) ;
END FUNC ;